`define hi

// comment

